/tech/tsmc/65LP/dig_libs/ARM_FEONLY/arm/tsmc/cln65lp/arm_tech/r2p0/lef/1p9m_6x2z/sc9_tech.lef