/project/tsmc65/shared/modified_libraries/tpdn65lpnv2od3_9lm.lef