//                          Copyright (C) 2015-2019 by EnICS Labs
//                      01
//                    01 10
//                   1 10 010101010              1010     0101010    1010101
//                   1 10         0              1  0    10     0   0      1
//                   1   1010101010              1  0   01  01010  1   10101
//                    010                        1  0   0  10      1  0
//                  01  01            01010101   1  0  1  01       1  01
//                 10 01 1010101010  10       0  1  0  1  0        10  10
//                 1  01          0  1   10   0  1  0  1  0         0    1
//                 10   01010101010  1  01 1  0  1  0  1  0          10   0
//                  01010            1  0  1  0  1  0  1  0           01   1
//                  0101             1  0  1  0  1  0  1  01           10  1
//                 1    0            1  0  1  0  1  0   0  10           0  1
//                0  10 01010101010  1  0  1  0  1  0   01  01010  10101   1
//                0 0 0           0  1  0  1  0  1  0    10     0  1      01
//                0 01  01010101010  1010  1010  1010     0101010  10101010
//                0    1
//                 1010
//                           ------<< System-on-Chip Lab >>-------
//
//       This module is confidential and proprietary property of EnICS Labs and the possession or use
//                      of this file requires a written license from EnICS Labs.


// ----------------------------------------------------------------------------------------------------------- 
// Project     : DVD_2019
// Title       : IO ring Verilog file for instantiation of the IO cells
// Filename    : ioring.v
// Author      : yuzhans
// Created     : December 29 2019 at 13:46:53
// ----------------------------------------------------------------------------------------------------------- 
// Description : Instantiation of all the required I/O cells.
// NOTE: This file generated by io_ring_xls_parse.py script applied on DVD_SoC_IOs.xlsx file
// ----------------------------------------------------------------------------------------------------------- 


module ioring (
                // Towards the package:
                PAD_CLOCK_EN,             // PAD #1
                PAD_TEST_EN,              // PAD #2
                PAD_IRAM_PROG_BYTE_0,     // PAD #6
                PAD_IRAM_PROG_BYTE_1,     // PAD #7
                PAD_IRAM_PROG_BYTE_2,     // PAD #8
                PAD_IRAM_PROG_BYTE_3,     // PAD #9
                PAD_IRAM_PROG_BYTE_4,     // PAD #10
                PAD_IRAM_PROG_BYTE_5,     // PAD #14
                PAD_IRAM_PROG_BYTE_6,     // PAD #15
                PAD_IRAM_PROG_BYTE_7,     // PAD #16
                PAD_FETCH_EN,             // PAD #17
                PAD_IRAM_PROG_BYTE_IDX_0, // PAD #18
                PAD_IRAM_PROG_BYTE_IDX_1, // PAD #22
                PAD_IRAM_PROG_DATA_BYTE,  // PAD #23
                PAD_CLK,                  // PAD #24
                PAD_RST_N,                // PAD #25
                PAD_DONE_FLAG,            // PAD #26
                PAD_IO_PLACEHOLD_30,      // PAD #30
                PAD_IO_PLACEHOLD_31,      // PAD #31
                PAD_IO_PLACEHOLD_32,      // PAD #32
                PAD_EXT_PERF_COUNTERS_5,  // PAD #33
                PAD_EXT_PERF_COUNTERS_6,  // PAD #34
                PAD_EXT_PERF_COUNTERS_0,  // PAD #38
                PAD_EXT_PERF_COUNTERS_1,  // PAD #39
                PAD_EXT_PERF_COUNTERS_2,  // PAD #40
                PAD_EXT_PERF_COUNTERS_3,  // PAD #41
                PAD_EXT_PERF_COUNTERS_4,  // PAD #42
                PAD_EXT_PERF_COUNTERS_7,  // PAD #46
                PAD_EXT_PERF_COUNTERS_8,  // PAD #47
                PAD_EXT_PERF_COUNTERS_9,  // PAD #48
                PAD_IO_PLACEHOLD_49,      // PAD #49
                PAD_IO_PLACEHOLD_50,      // PAD #50
                PAD_EXT_PERF_COUNTERS_10, // PAD #54
                PAD_EXT_PERF_COUNTERS_11, // PAD #55
                PAD_EXT_PERF_COUNTERS_12, // PAD #56
                PAD_EXT_PERF_COUNTERS_13, // PAD #57
                PAD_EXT_PERF_COUNTERS_14, // PAD #58
                PAD_EXT_PERF_COUNTERS_15, // PAD #62
                PAD_IRAM_PROG_WR,         // PAD #63
                PAD_IRAM_PROG_ADDR_BYTE,  // PAD #64

                // Towards the core:
                done_flag_from_core,
                clock_en_to_core,
                test_en_to_core,
                iram_prog_byte_to_core,
                fetch_en_to_core,
                iram_prog_byte_idx_to_core,
                iram_prog_data_byte_to_core,
                clk_to_core,
                rst_n_to_core,
                ext_perf_counters_to_core,
                iram_prog_wr_to_core,
                iram_prog_addr_byte_to_core
               );

   // External PADs toward the package:
   input  PAD_CLOCK_EN;             // PAD #1
   input  PAD_TEST_EN;              // PAD #2
   input  PAD_IRAM_PROG_BYTE_0;     // PAD #6
   input  PAD_IRAM_PROG_BYTE_1;     // PAD #7
   input  PAD_IRAM_PROG_BYTE_2;     // PAD #8
   input  PAD_IRAM_PROG_BYTE_3;     // PAD #9
   input  PAD_IRAM_PROG_BYTE_4;     // PAD #10
   input  PAD_IRAM_PROG_BYTE_5;     // PAD #14
   input  PAD_IRAM_PROG_BYTE_6;     // PAD #15
   input  PAD_IRAM_PROG_BYTE_7;     // PAD #16
   input  PAD_FETCH_EN;             // PAD #17
   input  PAD_IRAM_PROG_BYTE_IDX_0; // PAD #18
   input  PAD_IRAM_PROG_BYTE_IDX_1; // PAD #22
   input  PAD_IRAM_PROG_DATA_BYTE;  // PAD #23
   input  PAD_CLK;                  // PAD #24
   input  PAD_RST_N;                // PAD #25
   output PAD_DONE_FLAG;            // PAD #26
   output PAD_IO_PLACEHOLD_30;      // PAD #30
   output PAD_IO_PLACEHOLD_31;      // PAD #31
   output PAD_IO_PLACEHOLD_32;      // PAD #32
   input  PAD_EXT_PERF_COUNTERS_5;  // PAD #33
   input  PAD_EXT_PERF_COUNTERS_6;  // PAD #34
   input  PAD_EXT_PERF_COUNTERS_0;  // PAD #38
   input  PAD_EXT_PERF_COUNTERS_1;  // PAD #39
   input  PAD_EXT_PERF_COUNTERS_2;  // PAD #40
   input  PAD_EXT_PERF_COUNTERS_3;  // PAD #41
   input  PAD_EXT_PERF_COUNTERS_4;  // PAD #42
   input  PAD_EXT_PERF_COUNTERS_7;  // PAD #46
   input  PAD_EXT_PERF_COUNTERS_8;  // PAD #47
   input  PAD_EXT_PERF_COUNTERS_9;  // PAD #48
   output PAD_IO_PLACEHOLD_49;      // PAD #49
   output PAD_IO_PLACEHOLD_50;      // PAD #50
   input  PAD_EXT_PERF_COUNTERS_10; // PAD #54
   input  PAD_EXT_PERF_COUNTERS_11; // PAD #55
   input  PAD_EXT_PERF_COUNTERS_12; // PAD #56
   input  PAD_EXT_PERF_COUNTERS_13; // PAD #57
   input  PAD_EXT_PERF_COUNTERS_14; // PAD #58
   input  PAD_EXT_PERF_COUNTERS_15; // PAD #62
   input  PAD_IRAM_PROG_WR;         // PAD #63
   input  PAD_IRAM_PROG_ADDR_BYTE;  // PAD #64

   // Internal ports towards the logic core:
   input  done_flag_from_core;
   output clock_en_to_core;
   output test_en_to_core;
   output [7:0] iram_prog_byte_to_core;
   output fetch_en_to_core;
   output [1:0] iram_prog_byte_idx_to_core;
   output iram_prog_data_byte_to_core;
   output clk_to_core;
   output rst_n_to_core;
   output [15:0] ext_perf_counters_to_core;
   output iram_prog_wr_to_core;
   output iram_prog_addr_byte_to_core;

   // Inout direction control signals:

   wire logic_0;
   wire logic_1;

   hs_tielow  i_TIE_LOW  (.GROUND_TAP (logic_0));
   hs_tiehigh i_TIE_HIGH (.POWER_TAP  (logic_1));

   // Instantiation of IOs:

   // (1) IO ring corners:
   PCORNER i_PCORNER_NW ();
   PCORNER i_PCORNER_SW ();
   PCORNER i_PCORNER_SE ();
   PCORNER i_PCORNER_NE ();

   // (2) Power IOs:
   PVSS3CDG     i_VSSIO_3    (); //PAD #3
   PVDD2POC     i_VDDIO_4    (); //PAD #4
   PVDD1CDG     i_VDDCORE_5  (); //PAD #5
   PVDD1CDG     i_VDDCORE_11 (); //PAD #11
   PVDD2CDG     i_VDDIO_12   (); //PAD #12
   PVSS3CDG     i_VSSIO_13   (); //PAD #13
   PVSS3CDG     i_VSSIO_19   (); //PAD #19
   PVDD2CDG     i_VDDIO_20   (); //PAD #20
   PVDD1CDG     i_VDDCORE_21 (); //PAD #21
   PVSS3CDG     i_VSSIO_27   (); //PAD #27
   PVDD2CDG     i_VDDIO_28   (); //PAD #28
   PVDD1CDG     i_VDDCORE_29 (); //PAD #29
   PVSS3CDG     i_VSSIO_35   (); //PAD #35
   PVDD2CDG     i_VDDIO_36   (); //PAD #36
   PVDD1CDG     i_VDDCORE_37 (); //PAD #37
   PVSS3CDG     i_VSSIO_43   (); //PAD #43
   PVDD2CDG     i_VDDIO_44   (); //PAD #44
   PVDD1CDG     i_VDDCORE_45 (); //PAD #45
   PVSS3CDG     i_VSSIO_51   (); //PAD #51
   PVDD2CDG     i_VDDIO_52   (); //PAD #52
   PVDD1CDG     i_VDDCORE_53 (); //PAD #53
   PVSS3CDG     i_VSSIO_59   (); //PAD #59
   PVDD2CDG     i_VDDIO_60   (); //PAD #60
   PVDD1CDG     i_VDDCORE_61 (); //PAD #61

   // (3) Place-holder IOs:
   PDDW1216CDG  i_IO_PLACEHOLD_30 (.IE(logic_0), .C(), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_0), .PAD(PAD_IO_PLACEHOLD_30)); //PAD #30
   PDDW1216CDG  i_IO_PLACEHOLD_31 (.IE(logic_0), .C(), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_0), .PAD(PAD_IO_PLACEHOLD_31)); //PAD #31
   PDDW1216CDG  i_IO_PLACEHOLD_32 (.IE(logic_0), .C(), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_0), .PAD(PAD_IO_PLACEHOLD_32)); //PAD #32
   PDDW1216CDG  i_IO_PLACEHOLD_49 (.IE(logic_0), .C(), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_0), .PAD(PAD_IO_PLACEHOLD_49)); //PAD #49
   PDDW1216CDG  i_IO_PLACEHOLD_50 (.IE(logic_0), .C(), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_0), .PAD(PAD_IO_PLACEHOLD_50)); //PAD #50

   // (4) Digital IOs:

   //     [4.1] Inputs:
   PDDW1216SCDG i_CLOCK_EN             (.IE(logic_1), .C(clock_en_to_core             ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_CLOCK_EN            )); //PAD #1
   PDDW1216SCDG i_TEST_EN              (.IE(logic_1), .C(test_en_to_core              ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_TEST_EN             )); //PAD #2
   PDDW1216SCDG i_IRAM_PROG_BYTE_0     (.IE(logic_1), .C(iram_prog_byte_to_core[0]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_0    )); //PAD #6
   PDDW1216SCDG i_IRAM_PROG_BYTE_1     (.IE(logic_1), .C(iram_prog_byte_to_core[1]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_1    )); //PAD #7
   PDDW1216SCDG i_IRAM_PROG_BYTE_2     (.IE(logic_1), .C(iram_prog_byte_to_core[2]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_2    )); //PAD #8
   PDDW1216SCDG i_IRAM_PROG_BYTE_3     (.IE(logic_1), .C(iram_prog_byte_to_core[3]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_3    )); //PAD #9
   PDDW1216SCDG i_IRAM_PROG_BYTE_4     (.IE(logic_1), .C(iram_prog_byte_to_core[4]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_4    )); //PAD #10
   PDDW1216SCDG i_IRAM_PROG_BYTE_5     (.IE(logic_1), .C(iram_prog_byte_to_core[5]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_5    )); //PAD #14
   PDDW1216SCDG i_IRAM_PROG_BYTE_6     (.IE(logic_1), .C(iram_prog_byte_to_core[6]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_6    )); //PAD #15
   PDDW1216SCDG i_IRAM_PROG_BYTE_7     (.IE(logic_1), .C(iram_prog_byte_to_core[7]   ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_7    )); //PAD #16
   PDDW1216SCDG i_FETCH_EN             (.IE(logic_1), .C(fetch_en_to_core             ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_FETCH_EN            )); //PAD #17
   PDDW1216SCDG i_IRAM_PROG_BYTE_IDX_0 (.IE(logic_1), .C(iram_prog_byte_idx_to_core[0]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_IDX_0)); //PAD #18
   PDDW1216SCDG i_IRAM_PROG_BYTE_IDX_1 (.IE(logic_1), .C(iram_prog_byte_idx_to_core[1]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_BYTE_IDX_1)); //PAD #22
   PDDW1216SCDG i_IRAM_PROG_DATA_BYTE  (.IE(logic_1), .C(iram_prog_data_byte_to_core  ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_DATA_BYTE )); //PAD #23
   PDDW1216SCDG i_CLK                  (.IE(logic_1), .C(clk_to_core                  ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_CLK                 )); //PAD #24
   PDUW1216SCDG i_RST_N                (.IE(logic_1), .C(rst_n_to_core                ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_RST_N               )); //PAD #25
   PDDW1216SCDG i_EXT_PERF_COUNTERS_5  (.IE(logic_1), .C(ext_perf_counters_to_core[5]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_5 )); //PAD #33
   PDDW1216SCDG i_EXT_PERF_COUNTERS_6  (.IE(logic_1), .C(ext_perf_counters_to_core[6]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_6 )); //PAD #34
   PDDW1216SCDG i_EXT_PERF_COUNTERS_0  (.IE(logic_1), .C(ext_perf_counters_to_core[0]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_0 )); //PAD #38
   PDDW1216SCDG i_EXT_PERF_COUNTERS_1  (.IE(logic_1), .C(ext_perf_counters_to_core[1]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_1 )); //PAD #39
   PDDW1216SCDG i_EXT_PERF_COUNTERS_2  (.IE(logic_1), .C(ext_perf_counters_to_core[2]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_2 )); //PAD #40
   PDDW1216SCDG i_EXT_PERF_COUNTERS_3  (.IE(logic_1), .C(ext_perf_counters_to_core[3]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_3 )); //PAD #41
   PDDW1216SCDG i_EXT_PERF_COUNTERS_4  (.IE(logic_1), .C(ext_perf_counters_to_core[4]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_4 )); //PAD #42
   PDDW1216SCDG i_EXT_PERF_COUNTERS_7  (.IE(logic_1), .C(ext_perf_counters_to_core[7]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_7 )); //PAD #46
   PDDW1216SCDG i_EXT_PERF_COUNTERS_8  (.IE(logic_1), .C(ext_perf_counters_to_core[8]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_8 )); //PAD #47
   PDDW1216SCDG i_EXT_PERF_COUNTERS_9  (.IE(logic_1), .C(ext_perf_counters_to_core[9]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_9 )); //PAD #48
   PDDW1216SCDG i_EXT_PERF_COUNTERS_10 (.IE(logic_1), .C(ext_perf_counters_to_core[10]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_10)); //PAD #54
   PDDW1216SCDG i_EXT_PERF_COUNTERS_11 (.IE(logic_1), .C(ext_perf_counters_to_core[11]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_11)); //PAD #55
   PDDW1216SCDG i_EXT_PERF_COUNTERS_12 (.IE(logic_1), .C(ext_perf_counters_to_core[12]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_12)); //PAD #56
   PDDW1216SCDG i_EXT_PERF_COUNTERS_13 (.IE(logic_1), .C(ext_perf_counters_to_core[13]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_13)); //PAD #57
   PDDW1216SCDG i_EXT_PERF_COUNTERS_14 (.IE(logic_1), .C(ext_perf_counters_to_core[14]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_14)); //PAD #58
   PDDW1216SCDG i_EXT_PERF_COUNTERS_15 (.IE(logic_1), .C(ext_perf_counters_to_core[15]), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_EXT_PERF_COUNTERS_15)); //PAD #62
   PDDW1216SCDG i_IRAM_PROG_WR         (.IE(logic_1), .C(iram_prog_wr_to_core         ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_WR        )); //PAD #63
   PDDW1216SCDG i_IRAM_PROG_ADDR_BYTE  (.IE(logic_1), .C(iram_prog_addr_byte_to_core  ), .PE(logic_1), .DS(logic_1), .I(logic_0), .OEN(logic_1), .PAD(PAD_IRAM_PROG_ADDR_BYTE )); //PAD #64

   //     [4.2] Inouts: NONE

   //     [4.3] Outputs:
   PDUW1216SCDG i_DONE_FLAG (.IE(logic_0), .C( ), .PE(logic_1), .DS(logic_1), .I(done_flag_from_core ), .OEN(logic_0), .PAD(PAD_DONE_FLAG)); //PAD #26

endmodule

module hs_tielow (GROUND_TAP);
   output GROUND_TAP;
   assign GROUND_TAP = 1'b0;
endmodule

module hs_tiehigh (POWER_TAP);
   output POWER_TAP;
   assign POWER_TAP = 1'b1;
endmodule
